#include <stdio.h>

int print_stuff() {
    printf("Stuff\n");
    return 0;
}
